* Created by KLayout

* cell TOP
* pin A
* pin VDD
* pin Q
* pin VCC
.SUBCKT TOP 1 2 3 4
* net 1 A
* net 2 VDD
* net 3 Q
* net 4 VCC
* device instance $1 r90 *1 15.7,-13 PMOS
M$1 2 1 3 2 PMOS L=1U W=3.4U AS=9.52P AD=9.52P PS=12.4U PD=12.4U
* device instance $2 r270 *1 15.7,-39.5 NMOS
M$2 4 1 3 4 NMOS L=1U W=3.4U AS=9.52P AD=9.52P PS=12.4U PD=12.4U
.ENDS TOP
